-----------------------------------------------------------------
-- --
--* @name module_name_ --
--* @project --
--* @file module_name_.vhd --
--* @author _author_ --
--* @creation_date _date_ --
--* @revision_date  _date_  --
-- --
-----------------------------------------------------------------
-- Description:
--
--* @description 
--------------------------------------------------------------
--
-- Changelog:
--* @change _date_ _author_ => First version
--

library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
---- synthesis translate_off
--library unisim;
--use unisim.vcomponents.all;
---- synthesis translate_on

entity module_name_ is
  generic (

  );
  port (
    -- Clocks and Reset
    -- Signals
  );
end module_name_;

architecture implementation of module_name_  is
  ------------------------------------------------------------------------------------------ 
  --  Constants 
  ------------------------------------------------------------------------------------------ 

  ------------------------------------------------------------------------------------------ 
  --  Components
  ------------------------------------------------------------------------------------------ 

  ------------------------------------------------------------------------------------------ 
  --  Signals
  ------------------------------------------------------------------------------------------ 

begin
end architecture implementation;
