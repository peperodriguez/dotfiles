/////////////////////////////////////////////////////////////////
// 
//* @name module_name_ 
//* @project 
//* @file module_name_.sv 
//* @author _author_ 
//* @creation_date  _date_ 
//* @revision_date  _date_  
// 
/////////////////////////////////////////////////////////////////
// Description:
//
//* @description 
/////////////////////////////////////////////////////////////////
//
// Changelog:
//* @change _date_ _author_ => First version
//

// `include "YourIncludeFileHere.h"

module module_name_
  #(
    parameter _PAR_0 = _PAR_0_VALUE,
              _PAR_1 = _PAR_1_VALUE
  )
  (
    //Clocks and Resets
    //Input signals
    input _in_s_0,
    input _in_s_2,
    //Output signals
    output  _out_s_0,
    output  _out_s_1
  );

endmodule
